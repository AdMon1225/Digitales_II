`include "QoS.v"
`include "QoSSynth.v"
`include "probador.v"
`include "cmos_cells.v"

module testbench();

